interface intf;
  
  logic [7:0]add;
  logic [7:0]data_in;
  logic [7:0]data_out;
  logic we;
  logic clk;
  
endinterface
